-- intro_qsys_gpio_lcd_0.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity intro_qsys_gpio_lcd_0 is
	generic (
		N : natural := 8
	);
	port (
		Clk        : in    std_logic                    := '0';             --          clock.clk
		Address    : in    std_logic_vector(2 downto 0) := (others => '0'); -- avalon_slave_0.address
		ChipSelect : in    std_logic                    := '0';             --               .chipselect
		Read       : in    std_logic                    := '0';             --               .read
		Write      : in    std_logic                    := '0';             --               .write
		ReadData   : out   std_logic_vector(7 downto 0);                    --               .readdata
		WriteData  : in    std_logic_vector(7 downto 0) := (others => '0'); --               .writedata
		ParPort    : inout std_logic_vector(7 downto 0) := (others => '0'); --    conduit_end.export
		nReset     : in    std_logic                    := '0'              --     reset_sink.reset_n
	);
end entity intro_qsys_gpio_lcd_0;

architecture rtl of intro_qsys_gpio_lcd_0 is
	component ParallelPort is
		generic (
			N : natural := 8
		);
		port (
			Clk        : in    std_logic                    := 'X';             -- clk
			Address    : in    std_logic_vector(2 downto 0) := (others => 'X'); -- address
			ChipSelect : in    std_logic                    := 'X';             -- chipselect
			Read       : in    std_logic                    := 'X';             -- read
			Write      : in    std_logic                    := 'X';             -- write
			ReadData   : out   std_logic_vector(7 downto 0);                    -- readdata
			WriteData  : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			ParPort    : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			nReset     : in    std_logic                    := 'X'              -- reset_n
		);
	end component ParallelPort;

begin

	n_check : if N /= 8 generate
		assert false report "Supplied generics do not match expected generics" severity Failure;
	end generate;

	gpio_lcd_0 : component ParallelPort
		generic map (
			N => 8
		)
		port map (
			Clk        => Clk,        --          clock.clk
			Address    => Address,    -- avalon_slave_0.address
			ChipSelect => ChipSelect, --               .chipselect
			Read       => Read,       --               .read
			Write      => Write,      --               .write
			ReadData   => ReadData,   --               .readdata
			WriteData  => WriteData,  --               .writedata
			ParPort    => ParPort,    --    conduit_end.export
			nReset     => nReset      --     reset_sink.reset_n
		);

end architecture rtl; -- of intro_qsys_gpio_lcd_0
